module mem_shim (
    input             clk,
    input             rst_n,        // Soft reset (Watchdog) - resets FSM and FIFOs
    input             hard_rst_n,   // Hard reset (Power-on) - unused, same signal as rst_n in emu.sv

    // MPEG2 Core memory request FIFO (read side) — clocked on clk (mem_clk)
    input       [1:0] mem_req_rd_cmd,
    input      [21:0] mem_req_rd_addr,
    input      [63:0] mem_req_rd_dta,
    output reg        mem_req_rd_en,
    input             mem_req_rd_valid,

    // MPEG2 Core memory response FIFO (write side) — clocked on clk (mem_clk)
    output reg [63:0] mem_res_wr_dta,
    output reg        mem_res_wr_en,
    input             mem_res_wr_almost_full,

    // DDR3 Controller Interface (Avalon-MM 64-bit)
    output     [28:0] ddr3_addr,
    output      [7:0] ddr3_burstcnt,
    output            ddr3_read,
    output            ddr3_write,
    output     [63:0] ddr3_writedata,
    output      [7:0] ddr3_byteenable,
    input      [63:0] ddr3_readdata,
    input             ddr3_readdatavalid,
    input             ddr3_waitrequest,

    // Debug outputs
    output     [3:0]  debug_state,
    output      [1:0] debug_saved_cmd,
    output            debug_sdram_busy,
    output            debug_sdram_ack,
    output    [15:0]  debug_rd_count,
    output    [15:0]  debug_wr_count,
    output    [15:0]  debug_rsp_count,
    output    [15:0]  debug_read_pend_cycles
);

    // Command encoding (from mem_codes.v)
    localparam CMD_NOOP    = 2'd0;
    localparam CMD_REFRESH = 2'd1;
    localparam CMD_READ    = 2'd2;
    localparam CMD_WRITE   = 2'd3;

    // ADDR_ERR sentinel (MP@HL profile): generated by mem_addr.v on decoder startup flush.
    // Forwarding this to DDR3 causes permanent waitrequest. Filter it here.
    localparam ADDR_ERR = 22'h1EFFFF;

    // =========================================================================
    // DDR3 Avalon-MM outputs (combinational assigns from registered regs)
    // =========================================================================
    reg        ram_read;
    reg        ram_write;
    reg [28:0] ram_address;
    reg [63:0] ram_writedata;

    assign ddr3_read       = ram_read;
    assign ddr3_write      = ram_write;
    assign ddr3_addr       = ram_address;
    assign ddr3_writedata  = ram_writedata;
    assign ddr3_burstcnt   = 8'd1;
    assign ddr3_byteenable = 8'hFF;

    // =========================================================================
    // 2-State FSM + Skid Buffer
    // =========================================================================
    // state=0 (IDLE): Accept new FIFO commands
    // state=1 (WAIT): Wait for DDR3 bridge acceptance (!waitrequest)
    //
    // Address formula: {7'b0011000, addr[21:0]} = DENSE formula
    //   - bits[28:25] = 0011 = window 3 (HPS-mapped to 0x30000000)
    //   - bits[24:3]  = {3'b000, addr[18:0]} (8-byte stride per word address unit)
    //   - bits[2:0]   = addr[2:0]
    // This is the DENSE formula (fixes 24 MB TrustZone boundary crossing).
    //
    // ADDR_ERR (22'h1EFFFF) is dropped: writes are silently discarded,
    // reads return a synthetic 64'd0 response. This prevents DDR3 bus stall on
    // decoder pipeline flush at startup.

    reg state;

    // Skid buffer — captures the FIFO word that appears 1 cycle after rd_en is
    // deasserted (standard mode FIFO 1-cycle latency).
    reg        saved_valid;
    reg  [1:0] saved_cmd;
    reg [21:0] saved_addr;
    reg [63:0] saved_dta;

    always @(posedge clk) begin
        if (!rst_n) begin
            state          <= 0;
            ram_read       <= 0;
            ram_write      <= 0;
            ram_address    <= 0;
            ram_writedata  <= 0;
            mem_req_rd_en  <= 0;
            mem_res_wr_en  <= 0;
            mem_res_wr_dta <= 0;
            saved_valid    <= 0;
            saved_cmd      <= 0;
            saved_addr     <= 0;
            saved_dta      <= 0;
        end
        else begin
            // -----------------------------------------------------------------
            // Response Path (always active, independent of FSM state)
            // -----------------------------------------------------------------
            mem_res_wr_en <= ddr3_readdatavalid;
            if (ddr3_readdatavalid)
                mem_res_wr_dta <= ddr3_readdata;

            // -----------------------------------------------------------------
            // Command Path FSM
            // -----------------------------------------------------------------
            if (!state) begin
                // =============================================================
                // S_IDLE: Process next command (skid buffer has priority)
                // =============================================================
                if (saved_valid && !mem_res_wr_almost_full) begin
                    case (saved_cmd)
                        CMD_WRITE: begin
                            if (saved_addr == ADDR_ERR) begin
                                // Drop ADDR_ERR write — do not forward to DDR3
                                saved_valid   <= 0;
                                mem_req_rd_en <= !mem_res_wr_almost_full;
                            end else begin
                                ram_write     <= 1;
                                ram_address   <= {7'b0011000, saved_addr};
                                ram_writedata <= saved_dta;
                                state         <= 1;
                                saved_valid   <= 0;
                                mem_req_rd_en <= 0;
                            end
                        end
                        CMD_READ: begin
                            if (saved_addr == ADDR_ERR) begin
                                // Synthetic 0 response — do not forward to DDR3
                                mem_res_wr_dta <= 64'd0;
                                mem_res_wr_en  <= 1'b1;
                                saved_valid    <= 0;
                                mem_req_rd_en  <= !mem_res_wr_almost_full;
                            end else begin
                                ram_read      <= 1;
                                ram_address   <= {7'b0011000, saved_addr};
                                state         <= 1;
                                saved_valid   <= 0;
                                mem_req_rd_en <= 0;
                            end
                        end
                        default: begin
                            // NOOP/REFRESH: consume and resume flow
                            saved_valid   <= 0;
                            mem_req_rd_en <= !mem_res_wr_almost_full;
                        end
                    endcase
                end
                else if (mem_req_rd_valid && !mem_res_wr_almost_full) begin
                    case (mem_req_rd_cmd)
                        CMD_WRITE: begin
                            if (mem_req_rd_addr == ADDR_ERR) begin
                                // Drop ADDR_ERR write — keep flowing
                                mem_req_rd_en <= !mem_res_wr_almost_full;
                            end else begin
                                ram_write     <= 1;
                                ram_address   <= {7'b0011000, mem_req_rd_addr};
                                ram_writedata <= mem_req_rd_dta;
                                state         <= 1;
                                mem_req_rd_en <= 0;
                            end
                        end
                        CMD_READ: begin
                            if (mem_req_rd_addr == ADDR_ERR) begin
                                // Synthetic 0 response — keep flowing
                                mem_res_wr_dta <= 64'd0;
                                mem_res_wr_en  <= 1'b1;
                                mem_req_rd_en  <= !mem_res_wr_almost_full;
                            end else begin
                                ram_read      <= 1;
                                ram_address   <= {7'b0011000, mem_req_rd_addr};
                                state         <= 1;
                                mem_req_rd_en <= 0;
                            end
                        end
                        default: mem_req_rd_en <= !mem_res_wr_almost_full;
                    endcase
                end
                else begin
                    // No commands — keep asking
                    mem_req_rd_en <= !mem_res_wr_almost_full;
                end
            end
            else begin
                // =============================================================
                // S_WAIT: Hold ram_read/write until bridge accepts
                // =============================================================
                if (!ddr3_waitrequest) begin
                    ram_read      <= 0;
                    ram_write     <= 0;
                    state         <= 0;
                    mem_req_rd_en <= !mem_res_wr_almost_full;
                end

                // Skid buffer capture: FIFO outputs a word 1 cycle after rd_en
                // was deasserted (standard mode FIFO latency). Capture it here.
                if (mem_req_rd_valid && !saved_valid) begin
                    saved_valid <= 1;
                    saved_cmd   <= mem_req_rd_cmd;
                    saved_addr  <= mem_req_rd_addr;
                    saved_dta   <= mem_req_rd_dta;
                end
            end
        end
    end

    // =========================================================================
    // Debug counters
    // =========================================================================
    reg [15:0] rd_count;
    reg [15:0] wr_count;
    reg [15:0] rsp_count;

    wire rd_accepted = ddr3_read  && !ddr3_waitrequest;
    wire wr_accepted = ddr3_write && !ddr3_waitrequest;

    always @(posedge clk) begin
        if (!rst_n) begin
            rd_count  <= 0;
            wr_count  <= 0;
            rsp_count <= 0;
        end else begin
            if (rd_accepted)        rd_count  <= rd_count  + 1'd1;
            if (wr_accepted)        wr_count  <= wr_count  + 1'd1;
            if (ddr3_readdatavalid) rsp_count <= rsp_count + 1'd1;
        end
    end

    // =========================================================================
    // Debug telemetry
    // =========================================================================
    // debug_state = {cmd[1:0], saved_valid, state}
    //   M:0 = NOOP/IDLE    M:1 = NOOP/WAIT
    //   M:9 = READ/WAIT    M:D = WRITE/WAIT (no skid)
    //   M:F = WRITE/WAIT + skid occupied
    reg [1:0] debug_cmd;
    always @* begin
        if (ram_write)              debug_cmd = CMD_WRITE;
        else if (ram_read)          debug_cmd = CMD_READ;
        else if (saved_valid)       debug_cmd = saved_cmd;
        else if (mem_req_rd_valid)  debug_cmd = mem_req_rd_cmd;
        else                        debug_cmd = CMD_NOOP;
    end

    assign debug_state            = {debug_cmd[1:0], saved_valid, state};
    assign debug_saved_cmd        = saved_valid ? saved_cmd : CMD_NOOP;
    assign debug_sdram_busy       = ddr3_waitrequest;
    assign debug_sdram_ack        = rd_accepted | wr_accepted;
    assign debug_rd_count         = rd_count;
    assign debug_wr_count         = wr_count;
    assign debug_rsp_count        = rsp_count;
    assign debug_read_pend_cycles = 16'd0;

endmodule
