��m o d u l e   m e m _ s h i m   (  
         i n p u t                           c l k ,  
         i n p u t                           r s t _ n ,  
  
         / /   M P E G 2   C o r e   m e m o r y   r e q u e s t   F I F O   ( r e a d   s i d e )   �� �   c l o c k e d   o n   c l k   ( m e m _ c l k )  
         i n p u t               [ 1 : 0 ]   m e m _ r e q _ r d _ c m d ,  
         i n p u t             [ 2 1 : 0 ]   m e m _ r e q _ r d _ a d d r ,  
         i n p u t             [ 6 3 : 0 ]   m e m _ r e q _ r d _ d t a ,  
         o u t p u t   r e g                 m e m _ r e q _ r d _ e n ,  
         i n p u t                           m e m _ r e q _ r d _ v a l i d ,  
  
         / /   M P E G 2   C o r e   m e m o r y   r e s p o n s e   F I F O   ( w r i t e   s i d e )   �� �   c l o c k e d   o n   c l k   ( m e m _ c l k )  
         o u t p u t   r e g   [ 6 3 : 0 ]   m e m _ r e s _ w r _ d t a ,  
         o u t p u t   r e g                 m e m _ r e s _ w r _ e n ,  
         i n p u t                           m e m _ r e s _ w r _ a l m o s t _ f u l l ,  
  
         / /   D D R 3   C o n t r o l l e r   I n t e r f a c e   ( A v a l o n - M M   6 4 - b i t )  
         o u t p u t           [ 2 8 : 0 ]   d d r 3 _ a d d r ,  
         o u t p u t             [ 7 : 0 ]   d d r 3 _ b u r s t c n t ,  
         o u t p u t                         d d r 3 _ r e a d ,  
         o u t p u t                         d d r 3 _ w r i t e ,  
         o u t p u t           [ 6 3 : 0 ]   d d r 3 _ w r i t e d a t a ,  
         o u t p u t             [ 7 : 0 ]   d d r 3 _ b y t e e n a b l e ,  
         i n p u t             [ 6 3 : 0 ]   d d r 3 _ r e a d d a t a ,  
         i n p u t                           d d r 3 _ r e a d d a t a v a l i d ,  
         i n p u t                           d d r 3 _ w a i t r e q u e s t ,  
  
         / /   D e b u g   o u t p u t s  
         o u t p u t           [ 3 : 0 ]     d e b u g _ s t a t e ,  
         o u t p u t                         d e b u g _ s d r a m _ b u s y ,  
         o u t p u t                         d e b u g _ s d r a m _ a c k ,  
         o u t p u t         [ 1 5 : 0 ]     d e b u g _ r d _ c o u n t ,  
         o u t p u t         [ 1 5 : 0 ]     d e b u g _ w r _ c o u n t  
 ) ;  
  
         / /   C o m m a n d   e n c o d i n g   ( f r o m   m e m _ c o d e s . v )  
         l o c a l p a r a m   C M D _ N O O P         =   2 ' d 0 ;  
         l o c a l p a r a m   C M D _ R E F R E S H   =   2 ' d 1 ;  
         l o c a l p a r a m   C M D _ R E A D         =   2 ' d 2 ;  
         l o c a l p a r a m   C M D _ W R I T E       =   2 ' d 3 ;  
  
         / /   = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = =  
         / /   D D R 3   A v a l o n - M M   o u t p u t s  
         / /   = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = =  
         r e g                 r a m _ r e a d ;  
         r e g                 r a m _ w r i t e ;  
         r e g   [ 2 8 : 0 ]   r a m _ a d d r e s s ;  
         r e g   [ 6 3 : 0 ]   r a m _ w r i t e d a t a ;  
  
         a s s i g n   d d r 3 _ r e a d               =   r a m _ r e a d ;  
         a s s i g n   d d r 3 _ w r i t e             =   r a m _ w r i t e ;  
         a s s i g n   d d r 3 _ a d d r               =   r a m _ a d d r e s s ;  
         a s s i g n   d d r 3 _ w r i t e d a t a     =   r a m _ w r i t e d a t a ;  
         a s s i g n   d d r 3 _ b u r s t c n t       =   8 ' d 1 ;  
         a s s i g n   d d r 3 _ b y t e e n a b l e   =   8 ' h F F ;  
  
         / /   = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = =  
         / /   F S M  
         / /   = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = =  
         / /   s t a t e = 0   ( I D L E ) :   A c c e p t   n e w   F I F O   c o m m a n d s  
         / /   s t a t e = 1   ( W A I T ) :   W a i t   f o r   t r a n s a c t i o n   a c c e p t a n c e   ( ! w a i t r e q u e s t )  
  
         r e g   s t a t e ;  
  
         / /   S k i d   b u f f e r   t o   c a p t u r e   t h e   c o m m a n d   t h a t   e x i t s   t h e   F I F O    
         / /   o n e   c y c l e   a f t e r   w e   d e a s s e r t   m e m _ r e q _ r d _ e n .  
         r e g                 s a v e d _ v a l i d ;  
         r e g   [ 1 : 0 ]     s a v e d _ c m d ;  
         r e g   [ 2 1 : 0 ]   s a v e d _ a d d r ;  
         r e g   [ 6 3 : 0 ]   s a v e d _ d t a ;  
  
         a l w a y s   @ ( p o s e d g e   c l k )   b e g i n  
                 i f   ( ! r s t _ n )   b e g i n  
                         s t a t e                   < =   0 ;  
                         r a m _ r e a d             < =   0 ;  
                         r a m _ w r i t e           < =   0 ;  
                         r a m _ a d d r e s s       < =   0 ;  
                         r a m _ w r i t e d a t a   < =   0 ;  
                         m e m _ r e q _ r d _ e n   < =   0 ;  
                         m e m _ r e s _ w r _ e n   < =   0 ;  
                         m e m _ r e s _ w r _ d t a   < =   0 ;  
                         s a v e d _ v a l i d   < =   0 ;  
                         s a v e d _ c m d   < =   0 ;  
                         s a v e d _ a d d r   < =   0 ;  
                         s a v e d _ d t a   < =   0 ;  
                 e n d  
                 e l s e   b e g i n  
                         / /   - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - -  
                         / /   R e s p o n s e   P a t h   ( A l w a y s   A c t i v e )  
                         / /   - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - -  
                         m e m _ r e s _ w r _ e n   < =   d d r 3 _ r e a d d a t a v a l i d ;  
                         i f   ( d d r 3 _ r e a d d a t a v a l i d )  
                                 m e m _ r e s _ w r _ d t a   < =   d d r 3 _ r e a d d a t a ;  
  
                         / /   - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - -  
                         / /   C o m m a n d   P a t h  
                         / /   - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - - -  
                         i f   ( ! s t a t e )   b e g i n  
                                 / /   I D L E   S t a t e  
                                  
                                 / /   P r i o r i t y :   P r o c e s s   S a v e d   R e q u e s t   - >   N e w   R e q u e s t  
                                 i f   ( s a v e d _ v a l i d   & &   ! m e m _ r e s _ w r _ a l m o s t _ f u l l )   b e g i n  
                                         / /   P r o c e s s   S a v e d   R e q u e s t  
                                         c a s e   ( s a v e d _ c m d )  
                                                 C M D _ W R I T E :   b e g i n  
                                                         r a m _ w r i t e           < =   1 ;  
                                                         r a m _ a d d r e s s       < =   { 4 ' b 0 1 1 0 ,   2 ' b 0 0 ,   s a v e d _ a d d r ,   1 ' b 0 } ;  
                                                         r a m _ w r i t e d a t a   < =   s a v e d _ d t a ;  
                                                         s t a t e                   < =   1 ;           / /   G o   t o   W A I T  
                                                         s a v e d _ v a l i d       < =   0 ;           / /   C o n s u m e d  
                                                         m e m _ r e q _ r d _ e n   < =   0 ;           / /   E n s u r e   E N   s t a y s   l o w  
                                                 e n d  
                                                 C M D _ R E A D :   b e g i n  
                                                         r a m _ r e a d             < =   1 ;  
                                                         r a m _ a d d r e s s       < =   { 4 ' b 0 1 1 0 ,   2 ' b 0 0 ,   s a v e d _ a d d r ,   1 ' b 0 } ;  
                                                         s t a t e                   < =   1 ;           / /   G o   t o   W A I T  
                                                         s a v e d _ v a l i d       < =   0 ;           / /   C o n s u m e d  
                                                         m e m _ r e q _ r d _ e n   < =   0 ;           / /   E n s u r e   E N   s t a y s   l o w  
                                                 e n d  
                                                 d e f a u l t :   b e g i n  
                                                         / /   N O O P / R E F R E S H   f r o m   S k i d :   C o n s u m e d ,   s t a y   i n   I D L E  
                                                         s a v e d _ v a l i d       < =   0 ;  
                                                         / /   I m m e d i a t e l y   c h e c k   F I F O   o r   e n a b l e   f l o w  
                                                         m e m _ r e q _ r d _ e n   < =   ! m e m _ r e s _ w r _ a l m o s t _ f u l l ;  
                                                 e n d  
                                         e n d c a s e  
                                 e n d  
                                 e l s e   i f   ( m e m _ r e q _ r d _ v a l i d   & &   ! m e m _ r e s _ w r _ a l m o s t _ f u l l )   b e g i n  
                                         / /   P r o c e s s   N e w   F I F O   R e q u e s t  
                                         c a s e   ( m e m _ r e q _ r d _ c m d )  
                                                 C M D _ W R I T E :   b e g i n  
                                                         r a m _ w r i t e           < =   1 ;  
                                                         r a m _ a d d r e s s       < =   { 4 ' b 0 0 1 1 ,   m e m _ r e q _ r d _ a d d r ,   3 ' b 0 0 0 } ;  
                                                         r a m _ w r i t e d a t a   < =   m e m _ r e q _ r d _ d t a ;  
                                                         s t a t e                   < =   1 ;           / /   G o   t o   W A I T  
                                                         m e m _ r e q _ r d _ e n   < =   0 ;           / /   S t o p   p o p p i n g  
                                                 e n d  
                                                 C M D _ R E A D :   b e g i n  
                                                         r a m _ r e a d             < =   1 ;  
                                                         r a m _ a d d r e s s       < =   { 4 ' b 0 0 1 1 ,   m e m _ r e q _ r d _ a d d r ,   3 ' b 0 0 0 } ;  
                                                         s t a t e                   < =   1 ;           / /   G o   t o   W A I T  
                                                         m e m _ r e q _ r d _ e n   < =   0 ;           / /   S t o p   p o p p i n g  
                                                 e n d  
                                                 / /   I g n o r e   N O O P / R E F R E S H ,   k e e p   p o p p i n g  
                                                 d e f a u l t :   m e m _ r e q _ r d _ e n   < =   ! m e m _ r e s _ w r _ a l m o s t _ f u l l ;  
                                         e n d c a s e  
                                 e n d  
                                 e l s e   b e g i n  
                                         / /   N o   r e q u e s t s ,   m a i n t a i n   f l o w  
                                         m e m _ r e q _ r d _ e n   < =   ! m e m _ r e s _ w r _ a l m o s t _ f u l l ;  
                                 e n d  
                         e n d  
                         e l s e   b e g i n  
                                 / /   W A I T   S t a t e  
                                 i f   ( ! d d r 3 _ w a i t r e q u e s t )   b e g i n  
                                         / /   T r a n s a c t i o n   A c c e p t e d  
                                         r a m _ r e a d     < =   0 ;  
                                         r a m _ w r i t e   < =   0 ;  
                                         s t a t e           < =   0 ;   / /   B a c k   t o   I D L E  
                                          
                                         / /   R e s u m e   f l o w   c o n t r o l   ( l o o k   a h e a d   f o r   n e x t   c y c l e )  
                                         m e m _ r e q _ r d _ e n   < =   ! m e m _ r e s _ w r _ a l m o s t _ f u l l ;  
                                 e n d  
                                  
                                 / /   D A T A   L O S S   F I X :   C a p t u r e   S k i d   D a t a  
                                 / /   I f   w e   e n t e r e d   W A I T ,   m e m _ r e q _ r d _ e n   w a s   d e a s s e r t e d   i n   p r e v i o u s   c y c l e .  
                                 / /   B u t   F I F O   l a t e n c y   m e a n s   v a l i d   d a t a   m i g h t   a p p e a r   N O W   ( 1   c y c l e   l a t e ) .  
                                 / /   W e   M U S T   c a p t u r e   i t .  
                                 i f   ( m e m _ r e q _ r d _ v a l i d   & &   ! s a v e d _ v a l i d )   b e g i n  
                                         s a v e d _ v a l i d   < =   1 ;  
                                         s a v e d _ c m d       < =   m e m _ r e q _ r d _ c m d ;  
                                         s a v e d _ a d d r     < =   m e m _ r e q _ r d _ a d d r ;  
                                         s a v e d _ d t a       < =   m e m _ r e q _ r d _ d t a ;  
                                 e n d  
                                 / /   E l s e :   S t a y   i n   W A I T ,   h o l d i n g   r a m _ r e a d / w r i t e / a d d r / d a t a   s t a b l e  
                         e n d  
                 e n d  
         e n d  
  
         / /   = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = =  
         / /   D e b u g  
         / /   = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = = =  
         r e g   [ 1 5 : 0 ]   r d _ c o u n t ;  
         r e g   [ 1 5 : 0 ]   w r _ c o u n t ;  
  
         w i r e   r d _ a c c e p t e d   =   d d r 3 _ r e a d     & &   ! d d r 3 _ w a i t r e q u e s t ;  
         w i r e   w r _ a c c e p t e d   =   d d r 3 _ w r i t e   & &   ! d d r 3 _ w a i t r e q u e s t ;  
  
         a l w a y s   @ ( p o s e d g e   c l k )   b e g i n  
                 i f   ( ! r s t _ n )   b e g i n  
                         r d _ c o u n t   < =   0 ;  
                         w r _ c o u n t   < =   0 ;  
                 e n d   e l s e   b e g i n  
                         i f   ( r d _ a c c e p t e d )   r d _ c o u n t   < =   r d _ c o u n t   +   1 ' d 1 ;  
                         i f   ( w r _ a c c e p t e d )   w r _ c o u n t   < =   w r _ c o u n t   +   1 ' d 1 ;  
                 e n d  
         e n d  
  
         a s s i g n   d e b u g _ s t a t e             =   { 3 ' b 0 0 0 ,   s t a t e } ;  
         a s s i g n   d e b u g _ s d r a m _ b u s y   =   d d r 3 _ w a i t r e q u e s t ;  
         a s s i g n   d e b u g _ s d r a m _ a c k     =   r d _ a c c e p t e d   |   w r _ a c c e p t e d ;  
         a s s i g n   d e b u g _ r d _ c o u n t       =   r d _ c o u n t ;  
         a s s i g n   d e b u g _ w r _ c o u n t       =   w r _ c o u n t ;  
  
 e n d m o d u l e  
 